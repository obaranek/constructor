0
0 0 0 0  0 r h 
0 0 0 0  0 r h 
0 0 0 0  0 r h 
0 0 0 0  0 r h 
2 12 2 10 4 9 1 8 5 7 3 2 4 4 1 5 1 8 0 11 2 9 0 6 3 11 2 3 3 4 4 10 1 6 0 3 0 5 
4
